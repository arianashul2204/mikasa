module and_gate(c,a,b);
    input a,b;
    output c;
    
    and g1(c,a,b);
    
endmodule