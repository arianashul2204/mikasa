module and_gate(c,a,b);
    input a,b;
    output c;
    
    assign c = a&b;
    
endmodule