module nor_gate(c,a,b);
    input a,b;
    output c;
    
    nor g1(c,a,b);
    
endmodule