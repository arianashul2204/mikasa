module not_gate(a,b);
input b;
output a;
assign a = !b;
endmodule