module not_gate(a,b);
input b;
output a;
not g1(a,b);
endmodule