module or_gate(c,a,b);
    input a,b;
    output c;
    
    or g1(c,a,b);
    
endmodule